`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/05/2017 04:19:48 AM
// Design Name: 
// Module Name: InvSubBytes
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InvSubBytes(
    x, y
    );
    input  [31:0] x;
    output [31:0] y;
    
    function [7:0] S;
    input    [7:0] x;
      case (x)
          0:S= 82;   1:S=  9;   2:S=106;   3:S=213;   4:S= 48;   5:S= 54;   6:S=165;   7:S= 56;
          8:S=191;   9:S= 64;  10:S=163;  11:S=158;  12:S=129;  13:S=243;  14:S=215;  15:S=251;
         16:S=124;  17:S=227;  18:S= 57;  19:S=130;  20:S=155;  21:S= 47;  22:S=255;  23:S=135;
         24:S= 52;  25:S=142;  26:S= 67;  27:S= 68;  28:S=196;  29:S=222;  30:S=233;  31:S=203;
         32:S= 84;  33:S=123;  34:S=148;  35:S= 50;  36:S=166;  37:S=194;  38:S= 35;  39:S= 61;
         40:S=238;  41:S= 76;  42:S=149;  43:S= 11;  44:S= 66;  45:S=250;  46:S=195;  47:S= 78;
         48:S=  8;  49:S= 46;  50:S=161;  51:S=102;  52:S= 40;  53:S=217;  54:S= 36;  55:S=178;
         56:S=118;  57:S= 91;  58:S=162;  59:S= 73;  60:S=109;  61:S=139;  62:S=209;  63:S= 37;
         64:S=114;  65:S=248;  66:S=246;  67:S=100;  68:S=134;  69:S=104;  70:S=152;  71:S= 22;
         72:S=212;  73:S=164;  74:S= 92;  75:S=204;  76:S= 93;  77:S=101;  78:S=182;  79:S=146;
         80:S=108;  81:S=112;  82:S= 72;  83:S= 80;  84:S=253;  85:S=237;  86:S=185;  87:S=218;
         88:S= 94;  89:S= 21;  90:S= 70;  91:S= 87;  92:S=167;  93:S=141;  94:S=157;  95:S=132;
         96:S=144;  97:S=216;  98:S=171;  99:S=  0; 100:S=140; 101:S=188; 102:S=211; 103:S= 10;
        104:S=247; 105:S=228; 106:S= 88; 107:S=  5; 108:S=184; 109:S=179; 110:S= 69; 111:S=  6;
        112:S=208; 113:S= 44; 114:S= 30; 115:S=143; 116:S=202; 117:S= 63; 118:S= 15; 119:S=  2;
        120:S=193; 121:S=175; 122:S=189; 123:S=  3; 124:S=  1; 125:S= 19; 126:S=138; 127:S=107;
        128:S= 58; 129:S=145; 130:S= 17; 131:S= 65; 132:S= 79; 133:S=103; 134:S=220; 135:S=234;
        136:S=151; 137:S=242; 138:S=207; 139:S=206; 140:S=240; 141:S=180; 142:S=230; 143:S=115;
        144:S=150; 145:S=172; 146:S=116; 147:S= 34; 148:S=231; 149:S=173; 150:S= 53; 151:S=133;
        152:S=226; 153:S=249; 154:S= 55; 155:S=232; 156:S= 28; 157:S=117; 158:S=223; 159:S=110;
        160:S= 71; 161:S=241; 162:S= 26; 163:S=113; 164:S= 29; 165:S= 41; 166:S=197; 167:S=137;
        168:S=111; 169:S=183; 170:S= 98; 171:S= 14; 172:S=170; 173:S= 24; 174:S=190; 175:S= 27;
        176:S=252; 177:S= 86; 178:S= 62; 179:S= 75; 180:S=198; 181:S=210; 182:S=121; 183:S= 32;
        184:S=154; 185:S=219; 186:S=192; 187:S=254; 188:S=120; 189:S=205; 190:S= 90; 191:S=244;
        192:S= 31; 193:S=221; 194:S=168; 195:S= 51; 196:S=136; 197:S=  7; 198:S=199; 199:S= 49;
        200:S=177; 201:S= 18; 202:S= 16; 203:S= 89; 204:S= 39; 205:S=128; 206:S=236; 207:S= 95;
        208:S= 96; 209:S= 81; 210:S=127; 211:S=169; 212:S= 25; 213:S=181; 214:S= 74; 215:S= 13;
        216:S= 45; 217:S=229; 218:S=122; 219:S=159; 220:S=147; 221:S=201; 222:S=156; 223:S=239;
        224:S=160; 225:S=224; 226:S= 59; 227:S= 77; 228:S=174; 229:S= 42; 230:S=245; 231:S=176;
        232:S=200; 233:S=235; 234:S=187; 235:S= 60; 236:S=131; 237:S= 83; 238:S=153; 239:S= 97;
        240:S= 23; 241:S= 43; 242:S=  4; 243:S=126; 244:S=186; 245:S=119; 246:S=214; 247:S= 38;
        248:S=225; 249:S=105; 250:S= 20; 251:S= 99; 252:S= 85; 253:S= 33; 254:S= 12; 255:S=125; 
      endcase
    endfunction
    
    assign y = {S(x[31:24]), S(x[23:16]), S(x[15: 8]), S(x[ 7: 0])};
endmodule
